mode calc_top(input logic clk,
)